library ieee;
use ieee.std_logic_1164.all;




-----	SUBBYTES STEP LUT
entity sbox_lut is 
	port(in_byte : in std_logic_vector(0 to 7);
		 out_byte : out std_logic_vector(0 to 7));
end sbox_lut;




architecture arc of sbox_lut is 
	begin 
		with in_byte select 
			out_byte <= "01100011" when "00000000",
						"01111100" when "00000001",
						"01110111" when "00000010",
						"01111011" when "00000011",
						"11110010" when "00000100",
						"01101011" when "00000101",
						"01101111" when "00000110",
						"11000101" when "00000111",
						"00110000" when "00001000",
						"00000001" when "00001001",
						"01100111" when "00001010",
						"00101011" when "00001011",
						"11111110" when "00001100",
						"11010111" when "00001101",
						"10101011" when "00001110",
						"01110110" when "00001111",
						"11001010" when "00010000",
						"10000010" when "00010001",
						"11001001" when "00010010",
						"01111101" when "00010011",
						"11111010" when "00010100",
						"01011001" when "00010101",
						"01000111" when "00010110",
						"11110000" when "00010111",
						"10101101" when "00011000",
						"11010100" when "00011001",
						"10100010" when "00011010",
						"10101111" when "00011011",
						"10011100" when "00011100",
						"10100100" when "00011101",
						"01110010" when "00011110",
						"11000000" when "00011111",
						"10110111" when "00100000",
						"11111101" when "00100001",
						"10010011" when "00100010",
						"00100110" when "00100011",
						"00110110" when "00100100",
						"00111111" when "00100101",
						"11110111" when "00100110",
						"11001100" when "00100111",
						"00110100" when "00101000",
						"10100101" when "00101001",
						"11100101" when "00101010",
						"11110001" when "00101011",
						"01110001" when "00101100",
						"11011000" when "00101101",
						"00110001" when "00101110",
						"00010101" when "00101111",
						"00000100" when "00110000",
						"11000111" when "00110001",
						"00100011" when "00110010",
						"11000011" when "00110011",
						"00011000" when "00110100",
						"10010110" when "00110101",
						"00000101" when "00110110",
						"10011010" when "00110111",
						"00000111" when "00111000",
						"00010010" when "00111001",
						"10000000" when "00111010",
						"11100010" when "00111011",
						"11101011" when "00111100",
						"00100111" when "00111101",
						"10110010" when "00111110",
						"01110101" when "00111111",
						"00001001" when "01000000",
						"10000011" when "01000001",
						"00101100" when "01000010",
						"00011010" when "01000011",
						"00011011" when "01000100",
						"01101110" when "01000101",
						"01011010" when "01000110",
						"10100000" when "01000111",
						"01010010" when "01001000",
						"00111011" when "01001001",
						"11010110" when "01001010",
						"10110011" when "01001011",
						"00101001" when "01001100",
						"11100011" when "01001101",
						"00101111" when "01001110",
						"10000100" when "01001111",
						"01010011" when "01010000",
						"11010001" when "01010001",
						"00000000" when "01010010",
						"11101101" when "01010011",
						"00100000" when "01010100",
						"11111100" when "01010101",
						"10110001" when "01010110",
						"01011011" when "01010111",
						"01101010" when "01011000",
						"11001011" when "01011001",
						"10111110" when "01011010",
						"00111001" when "01011011",
						"01001010" when "01011100",
						"01001100" when "01011101",
						"01011000" when "01011110",
						"11001111" when "01011111",
						"11010000" when "01100000",
						"11101111" when "01100001",
						"10101010" when "01100010",
						"11111011" when "01100011",
						"01000011" when "01100100",
						"01001101" when "01100101",
						"00110011" when "01100110",
						"10000101" when "01100111",
						"01000101" when "01101000",
						"11111001" when "01101001",
						"00000010" when "01101010",
						"01111111" when "01101011",
						"01010000" when "01101100",
						"00111100" when "01101101",
						"10011111" when "01101110",
						"10101000" when "01101111",
						"01010001" when "01110000",
						"10100011" when "01110001",
						"01000000" when "01110010",
						"10001111" when "01110011",
						"10010010" when "01110100",
						"10011101" when "01110101",
						"00111000" when "01110110",
						"11110101" when "01110111",
						"10111100" when "01111000",
						"10110110" when "01111001",
						"11011010" when "01111010",
						"00100001" when "01111011",
						"00010000" when "01111100",
						"11111111" when "01111101",
						"11110011" when "01111110",
						"11010010" when "01111111",
						"11001101" when "10000000",
						"00001100" when "10000001",
						"00010011" when "10000010",
						"11101100" when "10000011",
						"01011111" when "10000100",
						"10010111" when "10000101",
						"01000100" when "10000110",
						"00010111" when "10000111",
						"11000100" when "10001000",
						"10100111" when "10001001",
						"01111110" when "10001010",
						"00111101" when "10001011",
						"01100100" when "10001100",
						"01011101" when "10001101",
						"00011001" when "10001110",
						"01110011" when "10001111",
						"01100000" when "10010000",
						"10000001" when "10010001",
						"01001111" when "10010010",
						"11011100" when "10010011",
						"00100010" when "10010100",
						"00101010" when "10010101",
						"10010000" when "10010110",
						"10001000" when "10010111",
						"01000110" when "10011000",
						"11101110" when "10011001",
						"10111000" when "10011010",
						"00010100" when "10011011",
						"11011110" when "10011100",
						"01011110" when "10011101",
						"00001011" when "10011110",
						"11011011" when "10011111",
						"11100000" when "10100000",
						"00110010" when "10100001",
						"00111010" when "10100010",
						"00001010" when "10100011",
						"01001001" when "10100100",
						"00000110" when "10100101",
						"00100100" when "10100110",
						"01011100" when "10100111",
						"11000010" when "10101000",
						"11010011" when "10101001",
						"10101100" when "10101010",
						"01100010" when "10101011",
						"10010001" when "10101100",
						"10010101" when "10101101",
						"11100100" when "10101110",
						"01111001" when "10101111",
						"11100111" when "10110000",
						"11001000" when "10110001",
						"00110111" when "10110010",
						"01101101" when "10110011",
						"10001101" when "10110100",
						"11010101" when "10110101",
						"01001110" when "10110110",
						"10101001" when "10110111",
						"01101100" when "10111000",
						"01010110" when "10111001",
						"11110100" when "10111010",
						"11101010" when "10111011",
						"01100101" when "10111100",
						"01111010" when "10111101",
						"10101110" when "10111110",
						"00001000" when "10111111",
						"10111010" when "11000000",
						"01111000" when "11000001",
						"00100101" when "11000010",
						"00101110" when "11000011",
						"00011100" when "11000100",
						"10100110" when "11000101",
						"10110100" when "11000110",
						"11000110" when "11000111",
						"11101000" when "11001000",
						"11011101" when "11001001",
						"01110100" when "11001010",
						"00011111" when "11001011",
						"01001011" when "11001100",
						"10111101" when "11001101",
						"10001011" when "11001110",
						"10001010" when "11001111",
						"01110000" when "11010000",
						"00111110" when "11010001",
						"10110101" when "11010010",
						"01100110" when "11010011",
						"01001000" when "11010100",
						"00000011" when "11010101",
						"11110110" when "11010110",
						"00001110" when "11010111",
						"01100001" when "11011000",
						"00110101" when "11011001",
						"01010111" when "11011010",
						"10111001" when "11011011",
						"10000110" when "11011100",
						"11000001" when "11011101",
						"00011101" when "11011110",
						"10011110" when "11011111",
						"11100001" when "11100000",
						"11111000" when "11100001",
						"10011000" when "11100010",
						"00010001" when "11100011",
						"01101001" when "11100100",
						"11011001" when "11100101",
						"10001110" when "11100110",
						"10010100" when "11100111",
						"10011011" when "11101000",
						"00011110" when "11101001",
						"10000111" when "11101010",
						"11101001" when "11101011",
						"11001110" when "11101100",
						"01010101" when "11101101",
						"00101000" when "11101110",
						"11011111" when "11101111",
						"10001100" when "11110000",
						"10100001" when "11110001",
						"10001001" when "11110010",
						"00001101" when "11110011",
						"10111111" when "11110100",
						"11100110" when "11110101",
						"01000010" when "11110110",
						"01101000" when "11110111",
						"01000001" when "11111000",
						"10011001" when "11111001",
						"00101101" when "11111010",
						"00001111" when "11111011",
						"10110000" when "11111100",
						"01010100" when "11111101",
						"10111011" when "11111110",
						"00010110" when "11111111",
						UNAFFECTED when others;
end;